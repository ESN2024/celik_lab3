// celik_lab3_sys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module celik_lab3_sys (
		input  wire       clk_clk,                         //                      clk.clk
		output wire       key_irq_irq,                     //                  key_irq.irq
		input  wire       reset_reset_n,                   //                    reset.reset_n
		output wire [7:0] seg1_external_connection_export, // seg1_external_connection.export
		output wire [7:0] seg2_external_connection_export  // seg2_external_connection.export
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                            // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                         // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [17:0] nios2_gen2_0_data_master_address;                             // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                          // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                               // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                           // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [17:0] nios2_gen2_0_instruction_master_address;                      // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                         // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect;  // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_chipselect -> opencores_i2c_0:wb_stb_i
	wire   [7:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata;    // opencores_i2c_0:wb_dat_o -> mm_interconnect_0:opencores_i2c_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest; // opencores_i2c_0:wb_ack_o -> mm_interconnect_0:opencores_i2c_0_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address;     // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_address -> opencores_i2c_0:wb_adr_i
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write;       // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_write -> opencores_i2c_0:wb_we_i
	wire   [7:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata;   // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_writedata -> opencores_i2c_0:wb_dat_i
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;      // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;   // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram0_s1_chipselect;                         // mm_interconnect_0:RAM0_s1_chipselect -> RAM0:chipselect
	wire  [31:0] mm_interconnect_0_ram0_s1_readdata;                           // RAM0:readdata -> mm_interconnect_0:RAM0_s1_readdata
	wire  [13:0] mm_interconnect_0_ram0_s1_address;                            // mm_interconnect_0:RAM0_s1_address -> RAM0:address
	wire   [3:0] mm_interconnect_0_ram0_s1_byteenable;                         // mm_interconnect_0:RAM0_s1_byteenable -> RAM0:byteenable
	wire         mm_interconnect_0_ram0_s1_write;                              // mm_interconnect_0:RAM0_s1_write -> RAM0:write
	wire  [31:0] mm_interconnect_0_ram0_s1_writedata;                          // mm_interconnect_0:RAM0_s1_writedata -> RAM0:writedata
	wire         mm_interconnect_0_ram0_s1_clken;                              // mm_interconnect_0:RAM0_s1_clken -> RAM0:clken
	wire         mm_interconnect_0_seg2_s1_chipselect;                         // mm_interconnect_0:SEG2_s1_chipselect -> SEG2:chipselect
	wire  [31:0] mm_interconnect_0_seg2_s1_readdata;                           // SEG2:readdata -> mm_interconnect_0:SEG2_s1_readdata
	wire   [1:0] mm_interconnect_0_seg2_s1_address;                            // mm_interconnect_0:SEG2_s1_address -> SEG2:address
	wire         mm_interconnect_0_seg2_s1_write;                              // mm_interconnect_0:SEG2_s1_write -> SEG2:write_n
	wire  [31:0] mm_interconnect_0_seg2_s1_writedata;                          // mm_interconnect_0:SEG2_s1_writedata -> SEG2:writedata
	wire         mm_interconnect_0_seg1_s1_chipselect;                         // mm_interconnect_0:SEG1_s1_chipselect -> SEG1:chipselect
	wire  [31:0] mm_interconnect_0_seg1_s1_readdata;                           // SEG1:readdata -> mm_interconnect_0:SEG1_s1_readdata
	wire   [1:0] mm_interconnect_0_seg1_s1_address;                            // mm_interconnect_0:SEG1_s1_address -> SEG1:address
	wire         mm_interconnect_0_seg1_s1_write;                              // mm_interconnect_0:SEG1_s1_write -> SEG1:write_n
	wire  [31:0] mm_interconnect_0_seg1_s1_writedata;                          // mm_interconnect_0:SEG1_s1_writedata -> SEG1:writedata
	wire         mm_interconnect_0_key_s1_chipselect;                          // mm_interconnect_0:KEY_s1_chipselect -> KEY:chipselect
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                            // KEY:readdata -> mm_interconnect_0:KEY_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                             // mm_interconnect_0:KEY_s1_address -> KEY:address
	wire         mm_interconnect_0_key_s1_write;                               // mm_interconnect_0:KEY_s1_write -> KEY:write_n
	wire  [31:0] mm_interconnect_0_key_s1_writedata;                           // mm_interconnect_0:KEY_s1_writedata -> KEY:writedata
	wire         mm_interconnect_0_seg3_s1_chipselect;                         // mm_interconnect_0:SEG3_s1_chipselect -> SEG3:chipselect
	wire  [31:0] mm_interconnect_0_seg3_s1_readdata;                           // SEG3:readdata -> mm_interconnect_0:SEG3_s1_readdata
	wire   [1:0] mm_interconnect_0_seg3_s1_address;                            // mm_interconnect_0:SEG3_s1_address -> SEG3:address
	wire         mm_interconnect_0_seg3_s1_write;                              // mm_interconnect_0:SEG3_s1_write -> SEG3:write_n
	wire  [31:0] mm_interconnect_0_seg3_s1_writedata;                          // mm_interconnect_0:SEG3_s1_writedata -> SEG3:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                      // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                        // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                         // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                           // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                       // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         irq_mapper_receiver0_irq;                                     // opencores_i2c_0:wb_inta_o -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                     // timer_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                         // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [KEY:reset_n, SEG1:reset_n, SEG2:reset_n, SEG3:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, opencores_i2c_0:wb_rst_i, rst_translator:in_reset, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [RAM0:reset, mm_interconnect_0:RAM0_reset1_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                       // rst_controller_001:reset_req -> RAM0:reset_req
	wire         nios2_gen2_0_debug_reset_request_reset;                       // nios2_gen2_0:debug_reset_request -> rst_controller_001:reset_in1

	celik_lab3_sys_KEY key (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (),                                    // external_connection.export
		.irq        (key_irq_irq)                          //                 irq.irq
	);

	celik_lab3_sys_RAM0 ram0 (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_ram0_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_ram0_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_ram0_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_ram0_s1_write),        //       .write
		.readdata   (mm_interconnect_0_ram0_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_ram0_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_ram0_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	celik_lab3_sys_SEG1 seg1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_seg1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg1_s1_readdata),   //                    .readdata
		.out_port   (seg1_external_connection_export)       // external_connection.export
	);

	celik_lab3_sys_SEG1 seg2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_seg2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg2_s1_readdata),   //                    .readdata
		.out_port   (seg2_external_connection_export)       // external_connection.export
	);

	celik_lab3_sys_SEG1 seg3 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_seg3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg3_s1_readdata),   //                    .readdata
		.out_port   ()                                      // external_connection.export
	);

	celik_lab3_sys_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	celik_lab3_sys_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	opencores_i2c opencores_i2c_0 (
		.wb_clk_i   (clk_clk),                                                      //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                               //      clock_reset.reset
		.scl_pad_io (),                                                             //         export_0.export
		.sda_pad_io (),                                                             //                 .export
		.wb_adr_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver0_irq)                                      // interrupt_sender.irq
	);

	celik_lab3_sys_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	celik_lab3_sys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                       //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.RAM0_reset1_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                            //        RAM0_reset1_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                              //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                          //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                           //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                                 //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                             //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                                //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                            //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                          //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                       //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                   //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                          //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                      //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),       //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),         //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),          //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),      //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),     //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),   //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),    //                                         .chipselect
		.KEY_s1_address                                 (mm_interconnect_0_key_s1_address),                              //                                   KEY_s1.address
		.KEY_s1_write                                   (mm_interconnect_0_key_s1_write),                                //                                         .write
		.KEY_s1_readdata                                (mm_interconnect_0_key_s1_readdata),                             //                                         .readdata
		.KEY_s1_writedata                               (mm_interconnect_0_key_s1_writedata),                            //                                         .writedata
		.KEY_s1_chipselect                              (mm_interconnect_0_key_s1_chipselect),                           //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),        //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),          //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),           //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),       //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),      //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),     //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),    //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),    //                                         .debugaccess
		.opencores_i2c_0_avalon_slave_0_address         (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address),      //           opencores_i2c_0_avalon_slave_0.address
		.opencores_i2c_0_avalon_slave_0_write           (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write),        //                                         .write
		.opencores_i2c_0_avalon_slave_0_readdata        (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata),     //                                         .readdata
		.opencores_i2c_0_avalon_slave_0_writedata       (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata),    //                                         .writedata
		.opencores_i2c_0_avalon_slave_0_waitrequest     (~mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest), //                                         .waitrequest
		.opencores_i2c_0_avalon_slave_0_chipselect      (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect),   //                                         .chipselect
		.RAM0_s1_address                                (mm_interconnect_0_ram0_s1_address),                             //                                  RAM0_s1.address
		.RAM0_s1_write                                  (mm_interconnect_0_ram0_s1_write),                               //                                         .write
		.RAM0_s1_readdata                               (mm_interconnect_0_ram0_s1_readdata),                            //                                         .readdata
		.RAM0_s1_writedata                              (mm_interconnect_0_ram0_s1_writedata),                           //                                         .writedata
		.RAM0_s1_byteenable                             (mm_interconnect_0_ram0_s1_byteenable),                          //                                         .byteenable
		.RAM0_s1_chipselect                             (mm_interconnect_0_ram0_s1_chipselect),                          //                                         .chipselect
		.RAM0_s1_clken                                  (mm_interconnect_0_ram0_s1_clken),                               //                                         .clken
		.SEG1_s1_address                                (mm_interconnect_0_seg1_s1_address),                             //                                  SEG1_s1.address
		.SEG1_s1_write                                  (mm_interconnect_0_seg1_s1_write),                               //                                         .write
		.SEG1_s1_readdata                               (mm_interconnect_0_seg1_s1_readdata),                            //                                         .readdata
		.SEG1_s1_writedata                              (mm_interconnect_0_seg1_s1_writedata),                           //                                         .writedata
		.SEG1_s1_chipselect                             (mm_interconnect_0_seg1_s1_chipselect),                          //                                         .chipselect
		.SEG2_s1_address                                (mm_interconnect_0_seg2_s1_address),                             //                                  SEG2_s1.address
		.SEG2_s1_write                                  (mm_interconnect_0_seg2_s1_write),                               //                                         .write
		.SEG2_s1_readdata                               (mm_interconnect_0_seg2_s1_readdata),                            //                                         .readdata
		.SEG2_s1_writedata                              (mm_interconnect_0_seg2_s1_writedata),                           //                                         .writedata
		.SEG2_s1_chipselect                             (mm_interconnect_0_seg2_s1_chipselect),                          //                                         .chipselect
		.SEG3_s1_address                                (mm_interconnect_0_seg3_s1_address),                             //                                  SEG3_s1.address
		.SEG3_s1_write                                  (mm_interconnect_0_seg3_s1_write),                               //                                         .write
		.SEG3_s1_readdata                               (mm_interconnect_0_seg3_s1_readdata),                            //                                         .readdata
		.SEG3_s1_writedata                              (mm_interconnect_0_seg3_s1_writedata),                           //                                         .writedata
		.SEG3_s1_chipselect                             (mm_interconnect_0_seg3_s1_chipselect),                          //                                         .chipselect
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                          //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                            //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                         //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                        //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect)                        //                                         .chipselect
	);

	celik_lab3_sys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
